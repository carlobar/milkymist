module LUT(a,b,sel,out);


input a;
input b;
input sel;
output out;	



/*
always @(a or b or sel) begin
	case(sel)
		1'b0: 
			out = a;
		1'b1:
			out = b;
	endcase
end
*/


LUT3 LUT3_mux (.O (out),
                         .I0 (sel),
                         .I1 (a),
                         .I2 (b));
defparam LUT3_mux.INIT = 8'he4; 


endmodule
